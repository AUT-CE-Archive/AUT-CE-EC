** Profile: "SCHEMATIC1-Sim"  [ E:\INSTALLATION ROOT\ORCAD 9.2\Projects\EC_Project_3_Part_5\ec_project_3_part_5-SCHEMATIC1-Sim.sim ] 

** Creating circuit file "ec_project_3_part_5-SCHEMATIC1-Sim.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of e:\installation root\orcad 9.2\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 1000 0.001 1
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\ec_project_3_part_5-SCHEMATIC1.net" 


.END
