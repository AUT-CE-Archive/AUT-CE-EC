** Profile: "SCHEMATIC1-Part_4"  [ E:\INSTALLATION ROOT\ORCAD 9.2\Projects\EC_Project_3_Part_4\ec_project_3_part_4-schematic1-part_4.sim ] 

** Creating circuit file "ec_project_3_part_4-schematic1-part_4.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of e:\installation root\orcad 9.2\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM R 1 15 1 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\ec_project_3_part_4-SCHEMATIC1.net" 


.END
