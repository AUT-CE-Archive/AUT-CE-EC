** Profile: "SCHEMATIC1-Part_4_3"  [ e:\installation root\orcad 9.2\projects\ec_project_3_part_4\ec_project_3_part_4-schematic1-part_4_3.sim ] 

** Creating circuit file "ec_project_3_part_4-schematic1-part_4_3.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of e:\installation root\orcad 9.2\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.STEP LIN PARAM R1 1 10 1 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\ec_project_3_part_4-SCHEMATIC1.net" 


.END
